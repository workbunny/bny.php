module compile

import base

pub fn run()!
{
	base.app_path()
	println("开发中...")
}
