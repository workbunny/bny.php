module files

import net.http
import json
import os
import base

// $if !macos {
import kingbes.libgo
// }

struct Http {
	url string = 'http://tool.kllxs.top/'
}

struct Res {
pub:
	code int
	msg  string
	data []struct {
	pub:
		name string
		ext  string
		type string
		size string
	}
}

/**
 * 获取文件列表
 *
 * @param string path 路径
 * @return !Res
 */
pub fn search(path string) !Res {
	text := http.get_text(Http{}.url + 'search?path=${path}')
	return json.decode(Res, text) or { panic('获取文件列表信息有误') }
}

/**
 * 获取php cli路径
 *
 * @return string
 */
pub fn path_php_cli() string {
	mut path := '/php'
	if os.user_os() == 'windows' {
		path += '/windows/x86_64/cli'
	} else if os.user_os() == 'linux' {
		path += '/linux/${base.get_machine()}/cli'
	}else {
		path += '/macos/${base.get_machine()}/cli'
	}
	return path
}

pub fn download_file(url string, path string) ! {
	// 判断系统是否为macos
	$if macos {
		res := os.execute('curl -fLsS -o "${path}" "${url}" &>/dev/null && echo 1 || echo 0')
		if res.output.trim_space() == '0' {
			panic('下载文件失败')
		}
	}$else{
		res := libgo.download_file(url, path)
		if res != '' {
			panic(res)
		}
	}
}

/**
 * 下载文件
 *
 * @param string path 路径
 * @param string file 文件名
 * @param string dir 目录
 * @return !void
 */
pub fn download(path string, file string, dir string) ! {
	url := Http{}.url + 'download?path=${path}&file=${file}'
	
	// vlang本身存在bug
	/* params := http.DownloaderParams{}
	// 下载文件
	resp := http.download_file_with_progress(url, base.path_add(dir, file), params)!
	return resp */
	
	// 判断系统是否为macos
	$if macos {
		res := os.execute('curl -fLsS -o "${base.path_add(dir, file)}" "${url}" &>/dev/null && echo 1 || echo 0')
		if res.output.trim_space() == '0' {
			panic('下载文件失败')
		}
	}$else{
		res := libgo.download_file(url, base.path_add(dir, file))
		if res != '' {
			panic(res)
		}
	}

}